module f_comparator_tb;


endmodule